module d7s(
    input en,
    input [3:0] x,
    output [6:0] y
);
    always_comb
        if(en)
            case (x)
            4'h0: y <= ~7'b0111111;
            4'h1: y <= ~7'b0000110;
            4'h2: y <= ~7'b1011011;
            4'h3: y <= ~7'b1001111;
            4'h4: y <= ~7'b1100110;
            4'h5: y <= ~7'b1101101;
            4'h6: y <= ~7'b1111101;
            4'h7: y <= ~7'b0100111;
            4'h8: y <= ~7'b1111111;
            4'h9: y <= ~7'b1101111;
            4'hA: y <= ~7'b1110111;
            4'hB: y <= ~7'b1111100;
            4'hC: y <= ~7'b0111001;
            4'hD: y <= ~7'b1011110;
            4'hE: y <= ~7'b1111001;
            4'hF: y <= ~7'b1110001;
            endcase
        else
            y <= ~7'd0;

endmodule
