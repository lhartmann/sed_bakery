module top(
	inout logic AUD_ADCDAT,
	inout logic AUD_ADCLRCK,
	inout logic AUD_BCLK,
	inout logic AUD_DACDAT,
	inout logic AUD_DACLRCK,
	inout logic AUD_XCK,
	inout logic CLOCK_27,
	inout logic CLOCK_50,
	inout logic DRAM_ADDR[11:0],
	inout logic DRAM_BA_0,
	inout logic DRAM_BA_1,
	inout logic DRAM_CAS_N,
	inout logic DRAM_CKE,
	inout logic DRAM_CLK,
	inout logic DRAM_CS_N,
	inout logic DRAM_DQ[15:0],
	inout logic DRAM_LDQM,
	inout logic DRAM_RAS_N,
	inout logic DRAM_UDQM,
	inout logic DRAM_WE_N,
	inout logic ENET_CLK,
	inout logic ENET_CMD,
	inout logic ENET_CS_N,
	inout logic ENET_DATA[15:0],
	inout logic ENET_INT,
	inout logic ENET_RD_N,
	inout logic ENET_RST_N,
	inout logic ENET_WR_N,
	inout logic EXT_CLOCK,
	inout logic FL_ADDR[21:0],
	inout logic FL_CE_N,
	inout logic FL_DQ[7:0],
	inout logic FL_OE_N,
	inout logic FL_RST_N,
	inout logic FL_WE_N,
	inout logic GPIO_0[35:0],
	inout logic GPIO_0[35],
	inout logic GPIO_1[35:0],
	inout logic HEX0[6:0],
	inout logic HEX1[6:0],
	inout logic HEX2[6:0],
	inout logic HEX3[6:0],
	inout logic HEX4[6:0],
	inout logic HEX5[6:0],
	inout logic HEX6[6:0],
	inout logic HEX7[6:0],
	inout logic I2C_SCLK,
	inout logic I2C_SDAT,
	inout logic IRDA_RXD,
	inout logic IRDA_TXD,
	inout logic KEY[3:0],
	inout logic LCD_BLON,
	inout logic LCD_DATA[7:0],
	inout logic LCD_EN,
	inout logic LCD_ON,
	inout logic LCD_RS,
	inout logic LCD_RW,
	inout logic LEDG[8:0],
	inout logic LEDR[17:0],
	inout logic OTG_ADDR[1:0],
	inout logic OTG_CS_N,
	inout logic OTG_DACK0_N,
	inout logic OTG_DACK1_N,
	inout logic OTG_DATA[15:0],
	inout logic OTG_DREQ0,
	inout logic OTG_DREQ1,
	inout logic OTG_FSPEED,
	inout logic OTG_INT0,
	inout logic OTG_INT1,
	inout logic OTG_LSPEED,
	inout logic OTG_RD_N,
	inout logic OTG_RST_N,
	inout logic OTG_WR_N,
	inout logic PS2_CLK,
	inout logic PS2_DAT,
	inout logic SD_CLK,
	inout logic SD_CMD,
	inout logic SD_DAT,
	inout logic SD_DAT3,
	inout logic SRAM_ADDR[17:0],
	inout logic SRAM_CE_N,
	inout logic SRAM_DQ[15:0],
	inout logic SRAM_LB_N,
	inout logic SRAM_OE_N,
	inout logic SRAM_UB_N,
	inout logic SRAM_WE_N,
	inout logic SW[17:0],
	inout logic TCK,
	inout logic TCS,
	inout logic TD_DATA[7:0],
	inout logic TD_HS,
	inout logic TDI,
	inout logic TDO,
	inout logic TD_RESET,
	inout logic TD_VS,
	inout logic UART_RXD,
	inout logic UART_TXD,
	inout logic VGA_B[9:0],
	inout logic VGA_BLANK,
	inout logic VGA_CLK,
	inout logic VGA_G[9:0],
	inout logic VGA_HS,
	inout logic VGA_R[9:0],
	inout logic VGA_SYNC,
	inout logic VGA_VS
);

endmodule
